`timescale 1ns / 1ps
`include "definitions.vh"

module adder(
    input [`WORD-1:0] a_in,
    input [`WORD-1:0] b_in,
    output [`WORD-1:0] add_out
    );
    
    assign add_out = a_in + b_in;
    
endmodule
