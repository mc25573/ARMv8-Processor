`timescale 1ns / 1ps
`define CYCLE 10
`define WORD  64
`define INSTR_LEN 32
`define DMEMFILE  "H:/ELC3338/Team8/CompOrg_Spring2018_S1_Team8/testfiles/ramData.data"
`define IMEMFILE  "H:/ELC3338/Team8/CompOrg_Spring2018_S1_Team8/testfiles/instrData.data"
`define RMEMFILE  "H:/ELC3338/Team8/CompOrg_Spring2018_S1_Team8/testfiles//regData.data"
