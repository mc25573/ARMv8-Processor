`timescale 1ns / 1ps
`include "definitions.vh"

module adder(
    input [`WORD-1:0] Ain,
    input [`WORD-1:0] Bin,
    output [`WORD-1:0] add_out
    );
    
    assign add_out = Ain + Bin;
    
endmodule
